`ifndef GRAPHICS_PARAMETERS
`define GRAPHICS_PARAMETERS

`define GRASS_PERCENTAGE 30 // 30% of screen is grass
`define STARTING_SPEED 1 // recommended: 1

`endif // GRAPHICS_PARAMETERS