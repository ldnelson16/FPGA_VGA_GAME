`ifndef CLOCKING_PARAMETERS
`define CLOCKING_PARAMETERS

`define INPUT_CLOCK_SPEED 50000000 // 50 Mhz
`define PLL_OUTPUT_CLOCK_SPEED 147140000 // 147.14 MHz
`define REFRESH_RATE 60
`define REFRESH_MAX (`INPUT_CLOCK_SPEED / `REFRESH_RATE)

`endif // CLOCKING_PARAMETERS