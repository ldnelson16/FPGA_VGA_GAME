`ifndef CLOCKING_PARAMETERS
`define CLOCKING_PARAMETERS

`define INPUT_CLOCK_SPEED 50000000;
`define REFRESH_RATE 60;
`define REFRESH_MAX (INPUT_CLOCK_SPEED / REFRESH_RATE);

`endif // CLOCKING_PARAMETERS